`define RX_FIFO  4'h0
`define TX_FIFO  4'h4
`define STAT_REG 4'h8
`define CTRL_REG 4'hC

