`define RESET_CMD 8'b1000_1110
`define START_CMD 8'b1000_1100
`define HALT_CMD  8'b1000_1010
`define READ_CMD  8'b1000_1000
`define WRITE_CMD 8'b1000_0110